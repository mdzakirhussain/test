* circuit of Transimpedance amplifier
vin n1 0 sin 0 2.5u 0.01k
M1000 n2 n1 0 0 nfet w=.07u l=.03u 
M1001 n2 n6 n4 n4 pfet w=.11u l=.03u 
R1 n1 n2 10k
vref n6 0 dc 0.7
R2 n5 n7 150k
L1 n4 n5 50p
vdd n7 0 dc 0.9
C0 n2 0 7.80f ic=0
C1 n1 0 15.59f ic=0
C2 n4 0 7.14f ic=0
C3 n6 0 3.71f ic=0
C4 n1 0 250f ic=0
.tran 1p 0.4u
.control
run
*plot v(n4)
plot v(n2)
.endc
.MODEL nfet NMOS LEVEL=3 PHI=0.700000 TOX=3.0600E-08 XJ=0.200000U TPG=1 
+ VTO=0.5666 DELTA=8.7630E-01 LD=9.0910E-10 KP=7.7684E-05 
+ UO=688.4 THETA=1.1640E-01 RSH=1.0310E+01 GAMMA=0.5904 
+ NSUB=1.3370E+16 NFS=5.9090E+11 VMAX=1.9740E+05 ETA=9.3470E-02 
+ KAPPA=2.1020E-01 CGDO=5.0000E-11 CGSO=5.0000E-11 
+ CGBO=3.1008E-10 CJ=2.7477E-04 MJ=5.5020E-01 CJSW=1.9263E-10 
+ MJSW=1.0000E-01 PB=9.9000E-01 

.MODEL pfet PMOS LEVEL=3 PHI=0.700000 TOX=3.0600E-08 XJ=0.200000U TPG=-1 
+ VTO=-0.7996 DELTA=2.4370E+00 LD=1.1000E-09 KP=1.8891E-05 
+ UO=167.4 THETA=9.5600E-02 RSH=1.0210E+01 GAMMA=0.3265 
+ NSUB=4.0890E+15 NFS=7.1500E+11 VMAX=1.2590E+05 ETA=8.2820E-02 
+ KAPPA=5.5040E+00 CGDO=5.0000E-11 CGSO=5.0000E-11 
+ CGBO=3.2338E-10 CJ=2.8023E-04 MJ=4.6284E-01 CJSW=2.1036E-10 
+ MJSW=1.2846E-01 PB=9.0211E-01

.end
