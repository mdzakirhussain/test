***************NG spice Tutorial****************
***************************************************
**************************************************
.include cmos_130nm.txt

**********Netlist*******
vdd net1 gnd 1.5
rd net1  vout 10k
vg vin gnd 0.6
*M1 Drain Gate Source Body
M1 vout vin gnd gnd NMOS w=1u L=130n

*********************************
***********Analysis*******
.control 
*op
*print @M1[id]
*print @M1[gm]
*print v(vout)

************DC Sweep********
dc vg 0 1.5 0.01
plot v(vout)
.endc
.end
